




`ifndef __PARAMETERS_simulation_VH__
`define __PARAMETERS_simulation_VH__ 1





/////////////////////////////////////////////////////////////////////////////////////////////////////////////// tb/simulator defines

`define SIMULATION_TYPE_BEHAVIOURAL 1
//`define SIMULATION_TYPE_POST_SYNTH_FUNCTIONAL 1
	// ^ pick one 

`define SIMULATION_FUNCTION_PERFORMED "sha"
`define SIMULATION_TEST_NAME "256_1bl_fixed_16_cells"

`define SHA256  (1)

//`define SHA256_1_BLOCK_FIXED_MESG_16_BLOCKS_16_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_32_BLOCKS_16_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_64_BLOCKS_16_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_128_BLOCKS_16_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_256_BLOCKS_16_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_512_BLOCKS_16_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_1024_BLOCKS_16_CELLS  (1)

//`define SHA256_1_BLOCK_FIXED_MESG_32_BLOCKS_32_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_64_BLOCKS_32_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_128_BLOCKS_32_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_256_BLOCKS_32_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_512_BLOCKS_32_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_1024_BLOCKS_32_CELLS  (1)

//`define SHA256_1_BLOCK_FIXED_MESG_64_BLOCKS_64_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_128_BLOCKS_64_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_256_BLOCKS_64_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_512_BLOCKS_64_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_1024_BLOCKS_64_CELLS  (1)

//`define SHA256_1_BLOCK_FIXED_MESG_128_BLOCKS_128_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_256_BLOCKS_128_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_512_BLOCKS_128_CELLS  (1)
//`define SHA256_1_BLOCK_FIXED_MESG_1024_BLOCKS_128_CELLS  (1)


//`define SHA256_1_BLOCK_FIXED_MESG_16_MESG_16_CELLS  (1)
//`define SHA256_2_BLOCK_FIXED_MESG_16_MESG_16_CELLS  (1)
//`define SHA256_4_BLOCK_FIXED_MESG_16_MESG_16_CELLS  (1)
//`define SHA256_8_BLOCK_FIXED_MESG_16_MESG_16_CELLS  (1)
//`define SHA256_16_BLOCK_FIXED_MESG_16_MESG_16_CELLS  (1)
//`define SHA256_32_BLOCK_FIXED_MESG_16_MESG_16_CELLS  (1)
//`define SHA256_64_BLOCK_FIXED_MESG_16_MESG_16_CELLS   (1)
//`define SHA256_128_BLOCK_FIXED_MESG_16_MESG_16_CELLS  (1)
//`define SHA256_256_BLOCK_FIXED_MESG_16_MESG_16_CELLS  (1)




`define SIMULATION_NR_LINES_DATA_OUT_READ (128) 
    // for IO; blocks tb natural $stop() if not set properly;
`define SIMULATION_NR_DATA_OUT_READ (`SIMULATION_NR_LINES_DATA_OUT_READ * `ARRAY_NR_CELLS)
// ^ comment if not known or desired 
// it is usually: (`SIMULATION_NR_LINES_DATA_OUT_READ * `ARRAY_NR_CELLS)



















